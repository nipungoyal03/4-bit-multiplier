magic
tech scmos
timestamp 1668249953
<< metal1 >>
rect -142 417 -128 724
rect -52 421 -38 720
rect 230 437 244 742
rect 420 457 438 766
rect 1798 682 1816 739
rect 1943 609 1957 737
rect 1451 599 1965 609
rect 1440 598 1965 599
rect 2266 518 2277 726
rect 1448 516 2280 518
rect 1460 507 2280 516
rect 2305 469 2314 727
rect 2313 461 2314 469
rect 974 459 1000 460
rect 974 457 1003 459
rect 420 456 1003 457
rect 230 435 249 437
rect 421 435 1003 456
rect -142 380 -129 417
rect -52 413 -37 421
rect -50 386 -37 413
rect 231 407 249 435
rect 974 434 1003 435
rect 231 402 247 407
rect -207 372 -129 380
rect -206 260 -194 372
rect -51 370 178 386
rect 231 385 898 402
rect 872 379 898 385
rect 168 294 178 370
rect 167 288 296 294
rect 168 287 178 288
rect 875 285 898 379
rect 984 395 1003 434
rect 1892 396 1899 397
rect 1249 395 1899 396
rect 984 376 1899 395
rect 984 375 1003 376
rect 1890 374 1899 376
rect 1892 297 1899 374
rect 875 270 1074 285
rect -206 249 -155 260
rect -205 248 -155 249
rect 120 204 157 210
rect -292 166 -229 167
rect -292 156 -161 166
rect -235 155 -161 156
rect 249 146 301 153
rect 841 121 850 198
rect 1631 194 1643 198
rect 1014 141 1080 152
rect 1634 109 1640 194
rect 1861 162 1898 168
rect 2455 145 2461 201
rect 118 58 314 66
rect 952 58 1129 66
rect 1730 61 1811 66
rect 290 53 301 58
rect 285 45 558 53
rect 1093 50 1106 58
rect 1800 53 1809 61
rect 1797 52 2167 53
rect 1081 42 1337 50
rect 1797 46 2161 52
rect 1633 43 1640 44
rect 1633 35 1634 43
rect 156 25 157 33
rect 156 -45 164 25
rect 841 -44 850 16
rect 1633 -29 1640 35
rect 2455 -20 2461 1
rect 2545 -17 2554 69
<< m2contact >>
rect 1798 663 1816 682
rect 1440 599 1451 609
rect 1448 507 1460 516
rect 2305 461 2313 469
rect 157 204 164 210
rect -303 156 -292 167
rect 239 145 249 153
rect 1002 141 1014 152
rect 841 111 850 121
rect 558 105 565 110
rect 1337 104 1343 110
rect 1853 162 1861 168
rect 2455 139 2461 145
rect 1634 103 1640 109
rect 2161 108 2167 113
rect 558 44 565 53
rect 1337 42 1343 50
rect 2161 46 2167 52
rect 1634 35 1640 43
rect 157 25 164 34
rect 841 16 850 26
rect 2455 1 2461 9
<< metal2 >>
rect -303 684 -292 686
rect -303 683 324 684
rect -303 682 1571 683
rect -303 667 1798 682
rect -303 167 -292 667
rect 324 666 1798 667
rect 1190 665 1798 666
rect 240 609 251 656
rect 240 599 1440 609
rect 240 401 251 599
rect 1448 516 1460 517
rect 1448 421 1460 507
rect 1853 469 1861 470
rect 1853 462 2305 469
rect 239 400 251 401
rect 1002 409 1469 421
rect 157 34 164 204
rect 239 153 250 400
rect 249 145 250 153
rect 1002 152 1014 409
rect 1853 168 1861 462
rect 558 53 565 105
rect 841 26 850 111
rect 1337 50 1343 104
rect 1634 43 1640 103
rect 2161 52 2167 108
rect 2455 9 2461 139
use half_adder  half_adder_0
timestamp 1668239862
transform 1 0 -147 0 1 180
box -17 -145 268 153
use full_adder  full_adder_0
timestamp 1667841856
transform 1 0 704 0 1 200
box -414 -164 248 147
use full_adder  full_adder_1
timestamp 1667841856
transform 1 0 1482 0 1 200
box -414 -164 248 147
use full_adder  full_adder_2
timestamp 1667841856
transform 1 0 2306 0 1 203
box -414 -164 248 147
<< labels >>
rlabel metal1 158 -34 158 -34 1 S0
rlabel metal1 845 -37 845 -37 1 S1
rlabel metal1 1635 -18 1635 -18 1 S2
rlabel metal1 2459 -15 2459 -15 1 S3
rlabel metal1 2549 -12 2549 -12 7 carry
rlabel metal1 -136 702 -136 702 1 b0
rlabel metal1 -44 699 -44 699 1 b1
rlabel metal1 233 717 233 717 1 b2
rlabel metal1 428 713 428 713 1 b3
rlabel metal1 1803 705 1803 705 1 a0
rlabel metal1 1947 713 1947 713 1 a1
rlabel metal1 2272 689 2272 689 1 a2
rlabel metal1 2308 687 2308 687 1 a3
<< end >>
