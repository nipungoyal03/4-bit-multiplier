magic
tech scmos
timestamp 1668239862
<< polysilicon >>
rect 113 81 116 82
rect 127 81 130 82
rect 220 0 223 1
rect 234 0 237 1
rect 16 -1 19 0
rect 30 -1 33 0
rect 108 -86 111 -85
rect 122 -86 125 -85
rect 219 -145 222 -144
rect 233 -145 236 -144
<< metal1 >>
rect -17 106 108 111
rect 141 107 169 111
rect -17 105 65 106
rect -17 28 -8 105
rect 64 97 108 102
rect 64 29 69 97
rect -17 24 11 28
rect 44 25 69 29
rect 161 30 169 107
rect 161 25 215 30
rect 248 25 268 29
rect -17 15 11 21
rect -17 -64 -12 15
rect 64 -56 71 25
rect 165 21 215 22
rect 164 17 215 21
rect 164 -55 169 17
rect 63 -61 64 -56
rect 71 -61 103 -56
rect 135 -61 169 -55
rect 153 -62 169 -61
rect -17 -69 103 -64
rect -17 -71 19 -69
rect -17 -75 -12 -71
rect 64 -115 71 -78
rect 64 -120 214 -115
rect 246 -119 266 -115
rect 169 -123 176 -120
rect 169 -129 214 -123
<< m2contact >>
rect 64 -61 71 -56
rect 64 -78 71 -73
<< metal2 >>
rect 64 -73 71 -61
use nand  nand_1
timestamp 1594232584
transform 1 0 121 0 1 123
box -24 -41 28 30
use nand  nand_0
timestamp 1594232584
transform 1 0 24 0 1 41
box -24 -41 28 30
use nand  nand_3
timestamp 1594232584
transform 1 0 228 0 1 42
box -24 -41 28 30
use nand  nand_2
timestamp 1594232584
transform 1 0 116 0 1 -44
box -24 -41 28 30
use nand  nand_4
timestamp 1594232584
transform 1 0 227 0 1 -103
box -24 -41 28 30
<< labels >>
rlabel metal1 263 26 263 26 7 sum
rlabel metal1 260 -117 260 -117 1 c_out
rlabel metal1 0 25 0 25 1 va
rlabel metal1 -8 18 -8 18 1 vb
<< end >>
