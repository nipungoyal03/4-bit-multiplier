magic
tech scmos
timestamp 1668279136
<< metal1 >>
rect 6016 1330 6021 1333
rect 551 1325 2740 1330
rect 2745 1325 4324 1330
rect 4329 1325 6059 1330
rect 292 1285 2531 1290
rect 2536 1285 4115 1290
rect 4120 1285 5815 1290
rect 5570 1252 5575 1262
rect 10 1247 2294 1252
rect 2299 1247 3878 1252
rect 3883 1247 5575 1252
rect 5326 1212 5331 1215
rect -362 1207 5346 1212
rect -378 1180 699 1184
rect -378 1113 -374 1180
rect -367 1105 -362 1140
rect -6 1119 -2 1180
rect -365 1068 -362 1105
rect 5 1080 10 1152
rect 276 1142 280 1180
rect 287 1102 292 1160
rect 535 1140 539 1180
rect 546 1102 551 1157
rect 2050 1079 2055 1207
rect -299 -4296 -294 1029
rect 73 939 78 1041
rect 355 943 360 1065
rect 614 964 619 1065
rect 2283 1057 2287 1059
rect 2039 1053 2897 1057
rect 830 969 848 1033
rect 73 934 162 939
rect 157 911 162 934
rect 258 938 360 943
rect 539 959 619 964
rect 157 906 169 911
rect 164 837 169 906
rect 258 844 263 938
rect 539 841 544 959
rect 723 951 848 969
rect 723 848 741 951
rect 2039 894 2043 1053
rect 2050 852 2055 978
rect 2283 904 2287 1053
rect 2294 863 2299 939
rect 2520 915 2524 1053
rect 2531 869 2536 983
rect 2729 910 2733 1053
rect 2740 869 2745 976
rect 459 -4291 467 1
rect 1144 -501 1153 27
rect 1144 -510 1665 -501
rect 1656 -1010 1665 -510
rect 1656 -1019 1753 -1010
rect 1744 -1165 1753 -1019
rect 1936 -1149 1943 36
rect 2758 -591 2764 34
rect 1839 -1156 1943 -1149
rect 2163 -597 2764 -591
rect 2163 -1165 2169 -597
rect 2848 -888 2857 54
rect 2370 -897 2857 -888
rect 2370 -1138 2379 -897
rect 3634 -927 3639 1207
rect 3623 -954 4506 -950
rect 3623 -1091 3627 -954
rect 3634 -1135 3639 -1040
rect 3867 -1095 3871 -954
rect 3878 -1124 3883 -1012
rect 4104 -1090 4108 -954
rect 4115 -1118 4120 -1028
rect 4313 -1082 4317 -954
rect 4324 -1118 4329 -1025
rect 2316 -1147 2379 -1138
rect 2117 -1171 2169 -1165
rect 2043 -4313 2051 -1974
rect 2728 -2531 2737 -1966
rect 3520 -2387 3527 -1955
rect 3520 -2394 3613 -2387
rect 2728 -2540 3459 -2531
rect 3450 -2903 3459 -2540
rect 3288 -2912 3459 -2903
rect 3288 -3128 3297 -2912
rect 3288 -3137 3440 -3128
rect 3606 -3135 3613 -2394
rect 4342 -2399 4348 -1951
rect 3288 -3148 3297 -3137
rect 3524 -3142 3613 -3135
rect 3893 -2405 4348 -2399
rect 3893 -3173 3899 -2405
rect 4432 -2753 4441 -1951
rect 4048 -2762 4441 -2753
rect 4048 -3128 4057 -2762
rect 5326 -2978 5331 1207
rect 5570 -2964 5575 1247
rect 5807 -2977 5812 1285
rect 6016 -2958 6021 1325
rect 5315 -2998 6191 -2994
rect 5315 -3073 5319 -2998
rect 5326 -3108 5331 -3054
rect 5559 -3064 5563 -2998
rect 5570 -3097 5575 -3023
rect 5796 -3070 5800 -2998
rect 5807 -3091 5812 -3030
rect 6005 -3058 6009 -2998
rect 6016 -3091 6021 -3022
rect 4012 -3137 4057 -3128
rect 3820 -3179 3899 -3173
rect 3735 -4342 3743 -3944
rect 4420 -4342 4429 -3953
rect 5212 -4383 5219 -3926
rect 6034 -4387 6040 -3927
rect 6124 -4379 6133 -3921
<< m2contact >>
rect 546 1325 551 1330
rect 2740 1325 2745 1330
rect 4324 1325 4329 1330
rect 287 1285 292 1290
rect 2531 1285 2536 1290
rect 4115 1285 4120 1290
rect 5 1247 10 1252
rect 2294 1247 2299 1252
rect 3878 1247 3883 1252
rect -367 1207 -362 1212
rect -367 1140 -362 1145
rect 5 1152 10 1157
rect 287 1160 292 1165
rect 546 1157 551 1162
rect 2050 1074 2055 1079
rect 2050 978 2055 983
rect 2294 939 2299 944
rect 2531 983 2536 988
rect 2740 976 2745 981
rect 3634 -932 3639 -927
rect 3634 -1040 3639 -1035
rect 3878 -1012 3883 -1007
rect 4115 -1028 4120 -1023
rect 4324 -1025 4329 -1020
rect 5570 -2969 5575 -2964
rect 5326 -2983 5331 -2978
rect 6016 -2963 6021 -2958
rect 5807 -2982 5812 -2977
rect 5326 -3054 5331 -3049
rect 5570 -3023 5575 -3018
rect 5807 -3030 5812 -3025
rect 6016 -3022 6021 -3017
<< metal2 >>
rect 2740 1330 2745 1331
rect -367 1145 -362 1207
rect 5 1157 10 1247
rect 287 1165 292 1285
rect 546 1162 551 1325
rect 2531 1290 2536 1291
rect 2050 983 2055 1074
rect 2294 944 2299 1247
rect 2531 988 2536 1285
rect 2740 981 2745 1325
rect 4115 1290 4120 1291
rect 3634 -1035 3639 -932
rect 3878 -1007 3883 1247
rect 4115 -1023 4120 1285
rect 4324 -1020 4329 1325
rect 5326 -3049 5331 -2983
rect 5570 -3018 5575 -2969
rect 5807 -3025 5812 -2982
rect 6016 -3017 6021 -2963
use and  and_0
timestamp 1668259600
transform 1 0 -335 0 1 1038
box -43 -9 96 76
use and  and_1
timestamp 1668259600
transform 1 0 37 0 1 1050
box -43 -9 96 76
use and  and_2
timestamp 1668259600
transform 1 0 319 0 1 1072
box -43 -9 96 76
use and  and_3
timestamp 1668259600
transform 1 0 578 0 1 1072
box -43 -9 96 76
use main-block  main-block_0
timestamp 1668260695
transform 1 0 0 0 1 0
box 0 0 2868 915
use main-block  main-block_1
timestamp 1668260695
transform 1 0 1584 0 1 -1987
box 0 0 2868 915
use main-block  main-block_2
timestamp 1668260695
transform 1 0 3276 0 1 -3960
box 0 0 2868 915
<< labels >>
rlabel metal1 -297 -4291 -296 -4289 1 p0
rlabel metal1 339 1182 339 1182 5 b0
rlabel metal1 2416 1055 2416 1055 1 b1
rlabel metal1 3876 -953 3876 -953 1 b2
rlabel metal1 5741 -2996 5741 -2996 1 b3
rlabel metal1 837 1013 837 1016 1 zero
rlabel metal1 463 -4274 463 -4274 1 p1
rlabel metal1 2047 -4294 2047 -4294 1 p2
rlabel metal1 3740 -4299 3740 -4299 1 p3
rlabel metal1 4424 -4296 4424 -4296 1 p4
rlabel metal1 5216 -4295 5216 -4295 1 p5
rlabel metal1 6037 -4285 6037 -4285 1 p6
rlabel metal1 6129 -4293 6129 -4293 1 p7
rlabel metal1 2834 1210 2834 1210 1 a0
rlabel metal1 2847 1250 2847 1250 1 a1
rlabel metal1 2837 1287 2837 1287 1 a2
rlabel metal1 2824 1328 2824 1328 5 a3
<< end >>
